module triple(
  input [3:0] a,
  output [5:0] result
);
  assign result = 3 * a;
endmodule
